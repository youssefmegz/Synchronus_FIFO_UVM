package shared_pkg;

bit test_finished ;
integer error_count ;
integer correct_count ;

int RD_EN_ON_DIST=30;
int WR_EN_ON_DIST=70;

parameter FIFO_WIDTH = 16;
parameter FIFO_DEPTH = 8;




endpackage